`timescale 1ns/1ps  // 시뮬레이션 시간 단위: 1ns, 정밀도: 1ps

//===========================================================
// 80비트 RCA(16비트 RCA × 5개) 모듈 테스트벤치
//===========================================================
module tb_rca16_80;

    //===============================
    // 입력 신호 정의 (자극용 reg)
    //===============================
    reg [79:0] A, B;   // 80비트 피연산자 A, B
    reg Cin;           // 초기 Carry 입력

    //===============================
    // 출력 신호 정의 (관찰용 wire)
    //===============================
    wire [79:0] Sum;   // 80비트 덧셈 결과
    wire Cout;         // 최종 캐리 출력 (MSB 이후 자리의 캐리)

    //===============================
    // 테스트 대상 DUT (rca16_80) 인스턴스화
    //===============================
    rca16_80 uut (
        .A(A),
        .B(B),
        .Cin(Cin),
        .Sum(Sum),
        .Cout(Cout)
    );

    //===============================
    // 테스트 시나리오 정의
    //===============================
    initial begin
        // 콘솔 출력 헤더
        $display("=================================================================================================================");
        $display("Time\t\t\t\tA\t\t\t\t\t\tB\t\t\t\t\t\tCin | Sum\t\t\t\t\t\t\t\t\tCout");
        $display("=================================================================================================================");

        //-------------------------------------------------------
        // 테스트 1: A = 0, B = 0, Cin = 0
        // → 기대 결과: Sum = 0, Cout = 0
        //-------------------------------------------------------
        A = 80'd0; B = 80'd0; Cin = 0;
        #10 $display("%0t\t%h\t%h\t%b | %h\t%b", $time, A, B, Cin, Sum, Cout);

        //-------------------------------------------------------
        // 테스트 2: A 최대값, B = 0, Cin = 0
        // → 기대 결과: Sum = A, Cout = 0
        //-------------------------------------------------------
        A = 80'hFFFFFFFFFFFFFFFFFFFF; B = 80'd0; Cin = 0;
        #10 $display("%0t\t%h\t%h\t%b | %h\t%b", $time, A, B, Cin, Sum, Cout);

        //-------------------------------------------------------
        // 테스트 3: A = 0, B 최대값, Cin = 0
        // → 기대 결과: Sum = B, Cout = 0
        //-------------------------------------------------------
        A = 80'd0; B = 80'hFFFFFFFFFFFFFFFFFFFF; Cin = 0;
        #10 $display("%0t\t%h\t%h\t%b | %h\t%b", $time, A, B, Cin, Sum, Cout);

        //-------------------------------------------------------
        // 테스트 4: A = 1, B = 1, Cin = 1
        // → 기대 결과: Sum = 3, 캐리 전파 확인
        //-------------------------------------------------------
        A = 80'd1; B = 80'd1; Cin = 1;
        #10 $display("%0t\t%h\t%h\t%b | %h\t%b", $time, A, B, Cin, Sum, Cout);

        //-------------------------------------------------------
        // 테스트 5: A = 2^79, B = 2^79, Cin = 0
        // → MSB 자리 오버플로우 확인 (Sum = 0, Cout = 1)
        //-------------------------------------------------------
        A = 80'h80000000000000000000; B = 80'h80000000000000000000; Cin = 0;
        #10 $display("%0t\t%h\t%h\t%b | %h\t%b", $time, A, B, Cin, Sum, Cout);

        //-------------------------------------------------------
        // 테스트 6: A = 중간값, B = 중간값
        // → 중간값 + 중간값 = Sum 오버플로우 확인
        //-------------------------------------------------------
        A = 80'h7FFFFFFFFFFFFFFFFFFF; B = 80'h7FFFFFFFFFFFFFFFFFFF; Cin = 0;
        #10 $display("%0t\t%h\t%h\t%b | %h\t%b", $time, A, B, Cin, Sum, Cout);

        //===============================
        // 시뮬레이션 종료
        //===============================
        $finish;
    end

endmodule
